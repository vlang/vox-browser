module html
